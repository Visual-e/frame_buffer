// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


`timescale 1ps / 1ps

// -------------------------------------------------------------------
// Dual clock FIFO. N bits wide. 5 addr lines.
//
// Originally generated by one of Gregg's toys. Modified for our
// needs. Share And Enjoy.
// -------------------------------------------------------------------

module alt_st_mlab_dcfifo_ack #(
    parameter DATA_WIDTH = 128,
    parameter READY_THRESHOLD = 14,
    parameter SIM_EMULATE = 1'b0
) 
(
    input din_clk,
    input din_sclr,
    input din_wreq,
    input [DATA_WIDTH-1:0] din,
    output reg din_ready,

    input dout_clk,
    input dout_sclr,
    input dout_rreq,
    output reg dout_valid,
    output [DATA_WIDTH-1:0] dout
);

///////////////////////////////
// resets

reg din_sclr_r = 1'b0 /* synthesis dont_merge */;
always @(posedge din_clk) begin
    din_sclr_r <= din_sclr;
end

reg dout_sclr_r = 1'b0 /* synthesis dont_merge */;
always @(posedge dout_clk) begin
    dout_sclr_r <= dout_sclr;
end

reg dout_sclr_val_r = 1'b0 /* synthesis dont_merge */;
always @(posedge dout_clk) begin
    dout_sclr_val_r <= dout_sclr;
end

///////////////////////////////
// underflow prevention
wire qual_rreq;
reg  empty;

assign qual_rreq = (dout_rreq | !dout_valid) & !empty;

///////////////////////////////
// write pointer

wire [4:0] din_wptr;
alt_hiconnect_cnt5ic wr_ctr (
    .clk(din_clk),
    .inc(din_wreq),
    .sclr(din_sclr_r),
    .dout(din_wptr)
);
defparam wr_ctr .SIM_EMULATE = SIM_EMULATE;

///////////////////////////////
// read pointer

wire [4:0] dout_lookahead_rptr;

alt_hiconnect_cnt5il lookahead_rd_ctr (
    .clk(dout_clk),
    .inc(qual_rreq),
    .sload(dout_sclr_r),
    .sload_data(5'b1),
    .dout(dout_lookahead_rptr)
);
defparam lookahead_rd_ctr .SIM_EMULATE = SIM_EMULATE;

///////////////////////////////
// storage

localparam MEM_WIDTH = (DATA_WIDTH % 20 == 0) ? DATA_WIDTH :
                                               (DATA_WIDTH / 20 + 1) * 20;
localparam RAM_BLOCKS = MEM_WIDTH / 20;

genvar i;

wire [MEM_WIDTH-1:0] sized_din;
wire [MEM_WIDTH-1:0] sized_dout;
wire [DATA_WIDTH-1:0] dout_w;
wire [4:0] waddr;
wire [4:0] dout_rptr;
wire [4:0] dout_next_rptr;

assign sized_din = din;
assign dout_w = sized_dout[DATA_WIDTH-1:0];

assign waddr = din_wptr;

generate for (i = 0; i < RAM_BLOCKS; i=i+1) begin : mem

    reg [4:0] waddr_m = 5'b0 /* synthesis dont_merge */;
    always @(posedge din_clk) waddr_m <= waddr;

    reg [19:0] wdata_m = 20'b0 /* synthesis dont_merge */;
    always @(posedge din_clk) wdata_m <= sized_din[(i+1)*20-1:i*20];

    reg [4:0] raddr_m = 5'b0 /* synthesis dont_merge */;
    always @(posedge dout_clk) begin
        if (dout_sclr_r) begin
            raddr_m <= 5'b0;
        end else begin
            raddr_m <= (qual_rreq) ? dout_lookahead_rptr : raddr_m;
        end
    end

    if (i == 0) begin
        assign dout_rptr = raddr_m;
        assign dout_next_rptr = (qual_rreq) ? dout_lookahead_rptr : raddr_m;
    end

    alt_hiconnect_mlab m (
        .wclk(din_clk),
        .wena(1'b1),
        .waddr_reg(waddr_m),
        .wdata_reg(wdata_m),
        .raddr(raddr_m),
        .rdata(sized_dout[(i+1)*20-1:i*20])
    );
    defparam m .WIDTH = 20;
    defparam m .ADDR_WIDTH = 5;
    defparam m .SIM_EMULATE = SIM_EMULATE;

end
endgenerate

///////////////////////////////////
// pointer cross domain exchange

wire [4:0] dout_xwptr;
wire [4:0] din_xrptr;

alt_hiconnect_gpx5 gx0 (
    .din_clk(din_clk),
    .din(din_wptr),
    .dout_clk(dout_clk),
    .dout(dout_xwptr)
);
defparam gx0 .SIM_EMULATE = SIM_EMULATE;

alt_hiconnect_gpx5 gx1 (
    .din_clk(dout_clk),
    .din(dout_rptr),
    .dout_clk(din_clk),
    .dout(din_xrptr)
);
defparam gx1 .SIM_EMULATE = SIM_EMULATE;

///////////////////////////////////
// compute used words

reg [4:0] rusedw = 5'b0;
reg [4:0] wusedw = 5'b0;

always @(posedge dout_clk) begin
    rusedw <= dout_xwptr - dout_rptr;
end

always @(posedge din_clk) begin
    wusedw <= din_wptr - din_xrptr;
end

///////////////////////////////
// compute almost full signal

always @(posedge din_clk) begin
    din_ready <= (wusedw < READY_THRESHOLD);
end

///////////////////////////////////
// compute empty

always @(posedge dout_clk) begin
    empty <= (dout_xwptr == dout_next_rptr);
end

///////////////////////////////
// compute valid signal

always @(posedge dout_clk) begin
    if (dout_sclr_val_r) 
        dout_valid <= 1'b0;
    else if (dout_rreq | !dout_valid) 
        dout_valid <= !empty;
end

///////////////////////////////
// output registers

reg [MEM_WIDTH-1:0] dout_r = {MEM_WIDTH{1'b0}};

generate for (i = 0; i < RAM_BLOCKS; i=i+1) begin : oreg

    always @(posedge dout_clk) begin
        if (dout_rreq | !dout_valid) dout_r[(i+1)*20-1:i*20] <= dout_w[(i+1)*20-1:i*20];
    end

end endgenerate

assign dout = dout_r[DATA_WIDTH-1:0];

endmodule

